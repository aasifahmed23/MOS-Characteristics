* CMOS Inverter
VDD 2 0 DC 1.8V
VIN 1 0 DC 0V
MN 3 1 0 0 NMOD W=360n L=180n
MP 3 1 2 2 PMOD W=1080n L=180n
.DC VIN 0 1.8V 0.025V
.MODEL NMOD NMOS(VTO=0.7 KP= 51u)
.MODEL PMOD PMOS(VTO=-0.7 KP= 17u)
.PROBE 
.END
 
